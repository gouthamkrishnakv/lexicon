// LEXICON: Generated file
// MODULE not
// Type: MODULE FILE

module not_mod(
    // port lists for the module
);
    // -- BODY OF MODULE

endmodule
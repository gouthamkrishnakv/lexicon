// LEXICON: Generated file
// MODULE not
// Type: TEST BENCH FILE

// TIMESCALE: <time_unit>/<time_precision>
`timescale 1ps/1ps

module not_tb;
    // -- ADD REGISTERS AND WIRES HERE

    initial begin
        $dumpfile("not.vcd");
        // use $dumpvars(level, variables ...) function for viewing its waveforms.

    end
    
endmodule